
module bluemax_platform (
	clk_clk,
	pio_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	pio_export;
	input		reset_reset_n;
endmodule
